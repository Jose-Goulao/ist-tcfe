CIRCUIT_T2_2

.options savecurrents


*********************************************
*	 	data import
*********************************************

.include ../doc/Dados_ngs-2.txt


*********************************************
*		 op & print
*********************************************

.control
op


echo "op_TAB2"

print i(vaux)
print i(h1)
print all
print v(n5,n2)
print v(n5,n8)

echo "op_END2"


*********************************************
*		    close
*********************************************

quit
.endc

.end

