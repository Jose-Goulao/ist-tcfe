CIRCUIT_T4

.options savecurrents


*********************************************
*	declaracion of components
*********************************************

.include valores.txt

Vcc vcc 0 12.0
Vin in 0 0 ac 1.0 sin(0 10m 1k)
Rin in in2 {rin_v}

* input coupling capacitor
Ci in2 base {ci_v}

* bias circuit
R1 vcc base {r1_v}
R2 base 0 {r2_v}

* gain stage
Q1 coll base emit BC547A
Rc vcc coll {rc_v}
Re emit 0 {re_v}

* bypass capacitor
Cb emit 0 {cb_v}


* output stage
Q2 0 coll emit2 BC557A
Rout emit2 vcc {rout_v}

* output coupling capacitor
Co emit2 out {co_v}

* load
RL out 0 {rl_v}


*********************************************
*	    	     setup
*********************************************

.op
.end

.control

set hcopypscolor=0
set color0=white
set color1=black
set color2=red
set color3=blue
set color4=violet
set color5=rgb:3/8/0
set color6=rgb:4/0/0


*********************************************
*	    	      op
*********************************************
op

echo "geral_TAB"

print v(coll)
print v(emit)
print v(emit2)
print v(emit2)-v(coll)
print v(coll)-v(base)
print v(coll)-v(emit)
print v(base)-v(emit)

echo "geral_END"


*********************************************
*	  	trans & plot
*********************************************
tran 1e-5 1e-2

plot v(coll)
hardcopy vocoll.eps vdb(coll)
hardcopy vo1.eps v(out)


*********************************************
*	        freq & plot
*********************************************
ac dec 10 10 100MEG

plot vdb(coll)
plot vp(coll)
hardcopy vo1f.eps vdb(coll)

plot vdb(out)
plot vp(out)
*hardcopy vo2f.eps vdb(out)


*---------------------
echo''

meas ac max MAX vdb(out) from=10 to=100MEG

let Vgain = abs(max)

let aux = max - 3 

hardcopy vo2f.eps vdb(out) max-3

meas ac LCOF WHEN vdb(out) = aux RISE=1
meas ac UCOF WHEN vdb(out) = aux CROSS=LAST

let Bandw = UCOF-LCOF

*---------------------
echo''

plot abs(v(in2)[40]/vin#branch[40]/(-1000))
let Zin = v(in2)[40]/vin#branch[40]/(-1000)
*let Zin = v(in2)[40]/(v(in)[40]-v(in2)[40])/100*1000

echo "INPUTimp_TAB"
print Zin 
echo "INPUTimp_END"

*---------------------
echo''

let Cost(resistor) = {rin_v} + {r1_v} + {r2_v} + {rc_v} + {re_v} + {rout_v} + {rl_v}
let Cost(capacitor) = {ci_v} + {cb_v} + {co_v}
let Cost(transistor) = 0.1*(2)
let Cost = Cost(resistor) + Cost(capacitor) + Cost(transistor)

let Merit = (Vgain*Bandw)/(Cost*LCOF)

*---------------------
echo''

echo "merit_TAB"

print Vgain
print Bandw
print Cost
print LCOF
echo ' ---------- & -------------------- '
print Merit

echo "merit_END"
echo ''


*********************************************
*		    close
*********************************************

quit
.endc


