CIRCUIT_T4_OUT

.options savecurrents

*********************************************
*	declaration of components
*********************************************
.include valores.txt


Vcc vcc 0 5.0
Vee vee 0 -5.0
Vin in 0 0

X1 0 inv_in vcc vee out uA741

R1 in inv_in 1000
R2 inv_in out 10000

* new source
Vn out 0 0 ac 1.0 sin(0 10m 1k)


*********************************************
*		     op
*********************************************
.op
.end

.control


*********************************************
*	        freq & imp
*********************************************
ac dec 10 10 100MEG


let Zout = -v(out)[40]/i(Vn)[40]

echo ''
echo "Outimp_TAB"
echo "Zout = $&Zout"
echo "Outimp_END"
echo ''


*********************************************
*		    close
*********************************************

quit
.endc


