CIRCUITO_T1

*********************************************
*	declaracao das componentes
*********************************************
*nome	entr	saida	valor

R1	N002	N003	1.00359089673
R2	N001	N002	2.04298963569
R3 	N004	N002	3.02503141993
R4 	0	N004	4.05647775356
R5 	N004	N005	3.07781188185
R6 	0	N006	2.01277040929
R7 	N008	N007	1.01993304256

Va	N003	0	5.11402517827
Id	N008	N005	1.03896393154

Vaux	N006	N007	0

G1	N005	N001	N002	N004	8.33526265782

H1	N004	N008	Vaux	7.23768458527


*********************************************
*		    setup
*********************************************

.model P2model NPN(Bf=200, CJE=12pF, CJC=2pF)
.control

set hcopypscolor=0
set color0=white
set color1=black
set color2=red
set color3=blue
set color4=violet
set color5=rgb:3/8/0
set color6=rgb:4/0/0


*********************************************
*		'corre' e mostra
*********************************************

op

echo ""
echo "+---------------------------------------------------+"
echo "|     VALORES DE VOLTAGENS E CURRENTES(#branch)     |"
echo "+---------------------------------------------------+"
echo ""
echo "op_TAB"
print all
echo "op_END"
echo ""
echo "______________________________________________________"
echo ""

echo "A currente em Ic é a mesma que passa em Vaux e em Vc (H1) e:"
print i(vaux)
 
echo ""
echo "A diferenca de potencial em Ib (G1) é a mesma em R3 e:"
print n004-n002

echo ""
echo "______________________________________________________"
echo ""


*********************************************
*		analise trans
*********************************************
*como este circuito nao varia com o tempo
*os valores no infinito são iguais aos iniciais

*primeiro valor é o passo e o ultimo o tempo final
*vão aparecer os valores iniciais

tran 1 2

hardcopy trans.ps v(n001) v(n005)
echo trans_FIG

*para ver um valor a variar no tempo,
*escrever print ... depois de tran ...

echo "______________________________________________________"
echo ""

*********************************************
*		analise ac
*********************************************

*ac dec <nº passos> <vlr minimo> <vlr maximo>
ac dec 10 1 100

*hardcopy ....
hardcopy acm.ps v(n001)  v(n005)
echo acm_FIG
hardcopy acp.ps v(n001)
echo acp_FIG 

hardcopy zim.ps abs(i(va))
echo zim_FIG

echo "______________________________________________________"
echo ""

*********************************************
*		encerrar
*********************************************

quit
.endc

.end
