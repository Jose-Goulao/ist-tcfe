CIRCUIT_T4_OUT

.options savecurrents

*********************************************
*	declaration of components
*********************************************
.include valores.txt


Vcc vcc 0 5.0
Vee vee 0 -5.0
Vin N1 0 0

X1 N2 inv_in vcc vee out uA741

C1 N1 inv_in 220n

R1 N2 0 1k
R2 N2 out 100k
R3 inv_in 0 10k

* new source
Vn out 0 0 ac 1.0 sin(0 10m 1k)



*********************************************
*		     op
*********************************************
.op
.end

.control


*********************************************
*	        freq & imp
*********************************************
ac dec 10 10 100MEG


let Zout = -v(out)[40]/i(Vn)[40]
let ReZout = Re(Zout)
let ImZout = Im(Zout)
let AbsZout = Abs(Zout)


echo ''
echo "Outimp_TAB"
echo "Zout = $&ReZout + $&ImZout j"
echo "Abs(Zout) = $&AbsZout"
echo "Outimp_END"
echo ''


*********************************************
*		    close
*********************************************

quit
.endc


