CIRCUIT_T1

.options savecurrents

*********************************************
*	declaracion of components
*********************************************
*nome	entr	saida	valor

R1	N2	N3	1.00359089673
R2	N1	N2	2.04298963569
R3 	N4	N2	3.02503141993
R4 	0	N4	4.05647775356
R5 	N4	N5	3.07781188185
R6 	0	N6	2.01277040929
R7 	N8	N7	1.01993304256

Va	N3	0	5.11402517827
Id	N8	N5	1.03896393154

Vaux	N6	N7	0

G1	N5	N1	N2	N4	7.23768458527
H1	N4	N8	Vaux	8.33526265782


*********************************************
*		'runs' & shows
*********************************************
.control

op

echo "op_TAB"

print i(vaux)
print i(h1)
print all
print v(n2,n4)
print v(n4,n8)

echo "op_END"



*********************************************
*		    close
*********************************************

quit
.endc

.end

