CIRCUIT_T3

.options savecurrents


*********************************************
*	declaracion of components
*********************************************
*nome	entr	saida	valor

*Source + Transformers

V1	N004	N001	dc 0 SIN(0 230 50 0 0 0)

*L1 N003 0 368m
*L2 N001 N004 300m
*K L1 L2 0.99999999999999

*Envelope Dectetor Circuit

D1	N001	N002 Default
D2	N004	N002 Default
D3	0	N001 Default
D4	0	N004 Default

C1	N002	0	10u


*Voltage Regulator Circuit

R1	P001	N002	1k

D5	P001	P002	Default
D6	P002	P003	Default
D7	P003	P004	Default
D8	P004	P005	Default
D9	P005	P006	Default
D10	P006	P007	Default
D11	P007	P008	Default
D12	P008	P009	Default
D13	P009	P010	Default
D14	P010	P011	Default
D15	P011	P012	Default
D16	P012	P013	Default
D17	P013	P014	Default
D18	P014	P015	Default
D19	P015	P016	Default
D20	P016	P017	Default
D21	P017	0	Default

.model Default D


*********************************************
*		 op & print
*********************************************

.control

set hcopypscolor=0
set color0=white
set color1=black
set color2=red
set color3=blue
set color4=violet
set color5=rgb:3/8/0
set color6=rgb:4/0/0


*********************************************
*	    trans & plot & table
*********************************************

tran 0.00017 50m 0

plot v(p001) 12
hardcopy trans-Vout_VR_all.eps v(p001) 12


*---------------------
*---------------------

tran 0.00017 205m 5m


plot v(n002)
hardcopy trans-Vout_ED.eps v(n002)

plot v(p001) 12
hardcopy trans-Vout_VR.eps v(p001) 12

plot v(p001)-12 0
hardcopy trans-Vout_(ac+dc).eps v(p001)-12 0

*---------------------
echo''

meas tran yavg AVG v(p001) from=10m to=210m
let Vout(AVG) = yavg

meas tran ymax MAX v(p001) from=10m to=210m
let Vout(MAX) = ymax

meas tran ymin MIN v(p001) from=10m to=210m
let Vout(MIN) = ymin

let Ripple(Vout) = Vout(MAX) - Vout(MIN)

*---------------------
echo''

let Cost(resistor) = 1
let Cost(capacitor) = 10
let Cost(diode) = 0.1*16
let Cost = Cost(resistor) + Cost(capacitor) + Cost(diode)


let Merit = 1/(Ripple(Vout) + (Vout(AVG)-12) + 1u)/(Cost)


*---------------------
echo''

echo "trans_TAB"

print Vout(AVG)
print Vout(MAX)
print Vout(MIN)
print Ripple(Vout)

echo "trans_END"

*---------------------
echo''

echo "cost_TAB"

print Cost(resistor)
print Cost(capacitor)
print Cost(diode)
print Cost
echo ' -------------------- & -------------------- '
print Merit

echo "cost_END"
echo ''


*********************************************
*		    close
*********************************************

quit
.endc

.end


