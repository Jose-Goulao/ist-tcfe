CIRCUIT_T2

.options savecurrents


*********************************************
*	 	data import
*********************************************

.include ../doc/Dados_ngs-1.txt


*********************************************
*		 op & print
*********************************************

.control
op


echo "op-1_TAB"

print i(vaux)
print i(h1)
print all
print v(n5,n2)
print v(n5,n8)
print v(n6,n8)

echo "op-1_END"


*********************************************
*		    close
*********************************************

quit
.endc

.end

